//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 07-Apr-2024  1.0.0  DWW  Initial creation
//
// 03-Mar-2025  1.1.0  DWW  No longer sending test packets!
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 1;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;
localparam RTL_TYPE      = 121475;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_DAY   = 3;
localparam VERSION_MONTH = 27;
localparam VERSION_YEAR  = 2025;
